library IEEE;
use IEEE.STD_LOGIC_1164.all;

--Entity
entity NOTGate is
	port( inport : in std_logic;
			outport: out std_logic);
end NOTGate;

--Achictecture
architecture Behavioral of NOTGate is
begin 

	outport <= not inport;
	
end Behavioral;